module not_gate1b(
    input a,
    output result
);
    assign result = ~a;
endmodule
